-- ============================================================================
-- 温度解码器测试台 (Temperature Decoder Testbench)
-- 功能：验证 temp_decoder 模块的正确性
-- 测试值：0000 1100 1000 1000 (对应 25.1°C)
-- ============================================================================
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_temp_decoder is
end tb_temp_decoder;

architecture Behavioral of tb_temp_decoder is

    -- ========================================================================
    -- 组件声明
    -- ========================================================================
    component temp_decoder is
        Port (
            clk         : in  STD_LOGIC;
            rst         : in  STD_LOGIC;
            temp_data   : in  STD_LOGIC_VECTOR(15 downto 0);
            bcd_tens    : out STD_LOGIC_VECTOR(3 downto 0);
            bcd_units   : out STD_LOGIC_VECTOR(3 downto 0);
            bcd_tenth   : out STD_LOGIC_VECTOR(3 downto 0)
        );
    end component;

    -- ========================================================================
    -- 信号定义
    -- ========================================================================
    signal clk        : STD_LOGIC := '0';
    signal rst        : STD_LOGIC := '0';
    signal temp_data  : STD_LOGIC_VECTOR(15 downto 0) := (others => '0');
    signal bcd_tens   : STD_LOGIC_VECTOR(3 downto 0);
    signal bcd_units  : STD_LOGIC_VECTOR(3 downto 0);
    signal bcd_tenth  : STD_LOGIC_VECTOR(3 downto 0);

    -- 时钟周期
    constant CLK_PERIOD : time := 10 ns;

begin

    -- ========================================================================
    -- 实例化被测模块
    -- ========================================================================
    UUT: temp_decoder
        port map (
            clk       => clk,
            rst       => rst,
            temp_data => temp_data,
            bcd_tens  => bcd_tens,
            bcd_units => bcd_units,
            bcd_tenth => bcd_tenth
        );

    -- ========================================================================
    -- 时钟生成
    -- ========================================================================
    clk_process: process
    begin
        clk <= '0';
        wait for CLK_PERIOD/2;
        clk <= '1';
        wait for CLK_PERIOD/2;
    end process;

    -- ========================================================================
    -- 测试激励
    -- ========================================================================
    stim_process: process
    begin
        -- 初始复位
        rst <= '1';
        wait for CLK_PERIOD * 5;
        rst <= '0';
        wait for CLK_PERIOD * 5;

        -- ====================================================================
        -- 测试1：25°C
        -- 13位值：0 0001 1001 0000 = 0x190
        -- 16位数据：0000 1100 1000 0000 = 0x0C80
        -- 整数部分 (bits 14-7): 0001 1001 = 25
        -- 小数部分 (bits 6-3):  0000 = 0
        -- 期望输出：tens=2, units=5, tenth=0
        -- ====================================================================
        temp_data <= "0000110010000000";  -- 0x0C80 = 25.0°C
        wait for CLK_PERIOD * 50;

        -- ====================================================================
        -- 测试2：25.5°C
        -- 13位值：0 0001 1001 1000 = 0x198
        -- 16位数据：0000 1100 1100 0000 = 0x0CC0
        -- 整数部分：25, 小数部分：1000 = 0.5
        -- 期望输出：tens=2, units=5, tenth=5
        -- ====================================================================
        temp_data <= "0000110011000000";  -- 0x0CC0 = 25.5°C
        wait for CLK_PERIOD * 50;

        -- ====================================================================
        -- 测试3：105°C
        -- 13位值：0 0110 1001 0000 = 0x690
        -- 16位数据：0011 0100 1000 0000 = 0x3480
        -- 整数部分：0110 1001 = 105
        -- 期望输出：tens=0, units=5, tenth=0 (只显示个位和十分位，百位不显示)
        -- ====================================================================
        temp_data <= "0011010010000000";  -- 0x3480 = 105°C
        wait for CLK_PERIOD * 50;

        -- ====================================================================
        -- 测试4：0.5°C
        -- 13位值：0 0000 0000 1000 = 0x008
        -- 16位数据：0000 0000 0100 0000 = 0x0040
        -- 整数部分：0, 小数部分：1000 = 0.5
        -- 期望输出：tens=0, units=0, tenth=5
        -- ====================================================================
        temp_data <= "0000000001000000";  -- 0x0040 = 0.5°C
        wait for CLK_PERIOD * 50;

        -- ====================================================================
        -- 测试5：99.9375°C (接近最大两位数)
        -- 13位值：0 0110 0011 1111 = 0x63F
        -- 16位数据：0011 0001 1111 1000 = 0x31F8
        -- 整数部分：0110 0011 = 99, 小数部分：1111 = 0.9375 ≈ 9
        -- 期望输出：tens=9, units=9, tenth=9
        -- ====================================================================
        temp_data <= "0011000111111000";  -- 0x31F8 = 99.9°C
        wait for CLK_PERIOD * 50;

        -- 完成测试，保持最后状态
        wait;
    end process;

end Behavioral;
