-- ============================================================================
-- BCD 到 7段数码管解码器 (BCD to 7-Segment Decoder)
-- 功能：将4位BCD码转换为7段数码管显示信号
-- 
-- 7段数码管段位定义（低电平有效，共阳极）：
--       a
--      ---
--   f |   | b
--      -g-
--   e |   | c
--      ---
--       d
--
-- seg(6 downto 0) = "gfedcba"
-- ============================================================================
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity bcd2seg is
    Port (
        bcd     : in  STD_LOGIC_VECTOR(3 downto 0);     -- 4位BCD输入 (0-9)
        seg     : out STD_LOGIC_VECTOR(6 downto 0)      -- 7段输出 "gfedcba" (低电平点亮)
    );
end bcd2seg;

architecture Behavioral of bcd2seg is
begin

    -- ========================================================================
    -- BCD 到 7段解码（共阳极，低电平点亮）
    -- seg = "gfedcba"
    -- ========================================================================
    with bcd select
        seg <=
            "1000000" when "0000",  -- 0: 显示 0 (a,b,c,d,e,f亮, g灭)
            "1111001" when "0001",  -- 1: 显示 1 (b,c亮)
            "0100100" when "0010",  -- 2: 显示 2 (a,b,d,e,g亮)
            "0110000" when "0011",  -- 3: 显示 3 (a,b,c,d,g亮)
            "0011001" when "0100",  -- 4: 显示 4 (b,c,f,g亮)
            "0010010" when "0101",  -- 5: 显示 5 (a,c,d,f,g亮)
            "0000010" when "0110",  -- 6: 显示 6 (a,c,d,e,f,g亮)
            "1111000" when "0111",  -- 7: 显示 7 (a,b,c亮)
            "0000000" when "1000",  -- 8: 显示 8 (全亮)
            "0010000" when "1001",  -- 9: 显示 9 (a,b,c,d,f,g亮)
            "1111111" when others;  -- 其他: 全灭

end Behavioral;
