-- ============================================================================
-- 度数符号显示模块 (Degree Symbol Display)
-- 功能：输出度数符号 "°" 的7段数码管显示信号
-- 
-- 7段数码管段位定义（低电平有效，共阳极）：
--       a
--      ---
--   f |   | b
--      -g-
--   e |   | c
--      ---
--       d
--
-- 度数符号 "°" 只点亮 a, b, f, g 四段
-- seg(6 downto 0) = "gfedcba"
-- ============================================================================
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity degree_symbol is
    Port (
        seg     : out STD_LOGIC_VECTOR(6 downto 0)      -- 7段输出 "gfedcba" (低电平点亮)
    );
end degree_symbol;

architecture Behavioral of degree_symbol is
begin

    -- ========================================================================
    -- 度数符号 "°" 显示
    -- 点亮段: a, b, f, g
    -- seg = "gfedcba" = "0011100" (g=0亮, f=0亮, e=1灭, d=1灭, c=1灭, b=0亮, a=0亮)
    -- ========================================================================
    seg <= "0011100";  -- 显示 °

end Behavioral;
