-- ============================================================================
-- 温度解码器测试台 (Temperature Decoder Testbench)
-- 功能：验证 temp_decoder 模块的正确性
-- 测试值：0000 1100 1000 1000 (对应 25.1°C)
-- ============================================================================
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_temp_decoder is
end tb_temp_decoder;

architecture Behavioral of tb_temp_decoder is

    -- ========================================================================
    -- 组件声明
    -- ========================================================================
    component temp_decoder is
        Port (
            clk         : in  STD_LOGIC;
            rst         : in  STD_LOGIC;
            temp_data   : in  STD_LOGIC_VECTOR(15 downto 0);
            bcd_tens    : out STD_LOGIC_VECTOR(3 downto 0);
            bcd_units   : out STD_LOGIC_VECTOR(3 downto 0);
            bcd_tenth   : out STD_LOGIC_VECTOR(3 downto 0)
        );
    end component;

    -- ========================================================================
    -- 信号定义
    -- ========================================================================
    signal clk        : STD_LOGIC := '0';
    signal rst        : STD_LOGIC := '0';
    signal temp_data  : STD_LOGIC_VECTOR(15 downto 0) := (others => '0');
    signal bcd_tens   : STD_LOGIC_VECTOR(3 downto 0);
    signal bcd_units  : STD_LOGIC_VECTOR(3 downto 0);
    signal bcd_tenth  : STD_LOGIC_VECTOR(3 downto 0);

    -- 时钟周期
    constant CLK_PERIOD : time := 10 ns;

begin

    -- ========================================================================
    -- 实例化被测模块
    -- ========================================================================
    UUT: temp_decoder
        port map (
            clk       => clk,
            rst       => rst,
            temp_data => temp_data,
            bcd_tens  => bcd_tens,
            bcd_units => bcd_units,
            bcd_tenth => bcd_tenth
        );

    -- ========================================================================
    -- 时钟生成
    -- ========================================================================
    clk_process: process
    begin
        clk <= '0';
        wait for CLK_PERIOD/2;
        clk <= '1';
        wait for CLK_PERIOD/2;
    end process;

    -- ========================================================================
    -- 测试激励
    -- ========================================================================
    stim_process: process
    begin
        -- 初始复位
        rst <= '1';
        wait for CLK_PERIOD * 5;
        rst <= '0';
        wait for CLK_PERIOD * 5;

        -- ====================================================================
        -- 测试1：25.1°C
        -- 二进制值：0000 1100 1000 1000
        -- 分析：
        --   整数部分 (bits 15-7): 0 0001 1001 = 25
        --   小数部分 (bits 6-3):  0001 = 0.0625 ≈ 0.1
        -- 期望输出：tens=2, units=5, tenth=1
        -- ====================================================================
        temp_data <= "0000110010001000";  -- 0x0C88
        wait for CLK_PERIOD * 50;  -- 等待 binary_bcd 转换完成

        -- ====================================================================
        -- 测试2：20.5°C
        -- 整数部分：20 = 0001 0100
        -- 小数部分：0.5 = 1000 (8 * 0.0625)
        -- 期望输出：tens=2, units=0, tenth=5
        -- ====================================================================
        temp_data <= "0000101001000000";  -- 20.5°C
        wait for CLK_PERIOD * 50;

        -- ====================================================================
        -- 测试3：30.0°C
        -- 整数部分：30 = 0001 1110
        -- 小数部分：0.0 = 0000
        -- 期望输出：tens=3, units=0, tenth=0
        -- ====================================================================
        temp_data <= "0000111100000000";  -- 30.0°C
        wait for CLK_PERIOD * 50;

        -- ====================================================================
        -- 测试4：0.5°C
        -- 期望输出：tens=0, units=0, tenth=5
        -- ====================================================================
        temp_data <= "0000000001000000";  -- 0.5°C
        wait for CLK_PERIOD * 50;

        -- ====================================================================
        -- 测试5：99.9°C (接近最大值)
        -- 期望输出：tens=9, units=9, tenth=9, sign=0
        -- ====================================================================
        temp_data <= "0011000111111000";  -- 99.9°C
        wait for CLK_PERIOD * 50;

        -- 完成测试，保持最后状态
        wait;
    end process;

end Behavioral;
